--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   17:22:51 02/13/2018
-- Design Name:   
-- Module Name:   C:/Users/gmpgreen/CENG450_Project/Shift_Right_TB.vhd
-- Project Name:  RegFile_ALU
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: Barrel_Shift_Right
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY Shift_Right_TB IS
END Shift_Right_TB;
 
ARCHITECTURE behavior OF Shift_Right_TB IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT Barrel_Shift_Right
    PORT(
         input : IN  std_logic_vector(15 downto 0);
         shift : IN  std_logic_vector(3 downto 0);
         output : OUT  std_logic_vector(15 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal input : std_logic_vector(15 downto 0) := (others => '0');
   signal shift : std_logic_vector(3 downto 0) := (others => '0');

 	--Outputs
   signal output : std_logic_vector(15 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Barrel_Shift_Right PORT MAP (
          input => input,
          shift => shift,
          output => output
        );
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 10 ns;	

      wait for clk_period*10;

      -- insert stimulus here
		input <= x"ABCD";
		shift <= x"4";
		wait for clk_period*3;
		input <= x"0ACC";
		shift <= x"8";
		wait for clk_period*3;
		input <= x"CA38";
		shift <= x"2";
		wait for clk_period*3;
	   input <= x"6F0F";
		shift <= x"1";
		wait for clk_period*3;
	   input <= x"A53C";
		shift <= x"F";
		
		wait;
   end process;

END;
